class axil_base_test extends uvm_test;

  `uvm_component_utils(axil_base_test)

  axil_env env;

  function new(string name = "", uvm_component parent = null);
    super.new(name, parent);
  endfunction

  virtual function void build_phase(uvm_phase phase);
    super.build_phase(phase);
    env = axil_env::type_id::create("env", this);
  endfunction

endclass
