typedef uvm_sequencer#(axil_wseq_item) axil_wsqr;
typedef uvm_sequencer#(axil_rseq_item) axil_rsqr;
