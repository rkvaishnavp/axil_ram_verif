typedef uvm_sequencer#(axil_rseq_item) axil_rsqr;
