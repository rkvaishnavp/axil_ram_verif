class axil_ragent extends uvm_agent;

  axil_rdrv rdrv;
  axil_rcov rcov;
  axil_rsqr rsqr;

  `uvm_component_utils(axil_ragent)

endclass
