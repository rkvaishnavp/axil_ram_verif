class axil_rcov extends uvm_subscriber #(axil_rseq_item);
    
endclass
