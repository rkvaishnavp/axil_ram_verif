package axil_pkg;

  import uvm_pkg::*;
  

endpackage
