typedef uvm_sequencer#(axil_wseq_item) axil_wsqr;
